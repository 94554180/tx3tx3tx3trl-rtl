package tx3tx3trl_pkg;
endpackage
